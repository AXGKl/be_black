/tmp/black/pkgs/vim-8.1.0390-py37_8/share/vim/vim81/tutor/tutor.sv